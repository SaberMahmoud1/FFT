package twiddle_pkg;
    parameter TWIDDLE_SIZE = 16; 
    // localparam logic signed [TWIDDLE_SIZE-1:0] TWIDDLE_REAL [0:15] = '{
    //     16'sd32767,              //wo
    //     16'sd32138,              //w1
    //     16'sd30274,              //w2
    //     16'sd27245,              //w3
    //     16'sd23170,              //w4
    //     16'sd18204,
    //     16'sd12539,              //w6
    //     16'sd6393,
    //     16'sd0,                  //w8
    //     -16'sd6393,
    //     -16'sd12539,
    //     -16'sd18204,
    //     -16'sd23170,
    //     -16'sd27245,
    //     -16'sd30274,
    //     -16'sd32138
    // };

    // localparam logic signed [TWIDDLE_SIZE-1:0] TWIDDLE_IMAG [0:15] = '{
    //     16'sd0, -16'sd6393, -16'sd12539, -16'sd18204,
    //     -16'sd23170, -16'sd27245, -16'sd30274, -16'sd32138,
    //     -16'sd32768, -16'sd32138, -16'sd30274, -16'sd27245,
    //     -16'sd23170, -16'sd18204, -16'sd12539, -16'sd6393
    // };


// localparam logic signed [15:0] TWIDDLE_REAL [0:15] = '{
//     16'b0000000100000000, //  +256 (1.0)
//     16'b0000000011111011, //  +251
//     16'b0000000011101100, //  +236
//     16'b0000000011010100, //  +212
//     16'b0000000010110101, //  +181
//     16'b0000000010001110, //  +142
//     16'b0000000001100001, //  +97
//     16'b0000000000110001, //  +49
//     16'b0000000000000000, //  0
//     16'b1111111111001110, //  -50
//     16'b1111111110011110, //  -98
//     16'b1111111101110001, //  -113
//     16'b1111111101001010, //  -150
//     16'b1111111100101011, //  -173
//     16'b1111111100010011, //  -189
//     16'b1111111100000100  //  -252
// };

//     localparam logic signed [15:0] TWIDDLE_IMAG [0:15] = '{
//     16'b0000000000000000, //    0
//     16'b1111111111001110, //  -50
//     16'b1111111110011110, //  -98
//     16'b1111111101110001, // -113
//     16'b1111111101001010, // -150
//     16'b1111111100101011, // -173
//     16'b1111111100010011, // -189
//     16'b1111111100000100, // -252
//     16'b1111111100000000, // -256
//     16'b1111111100000100, // -252
//     16'b1111111100010011, // -189
//     16'b1111111100101011, // -173
//     16'b1111111101001010, // -150
//     16'b1111111101110001, // -113
//     16'b1111111110011110, //  -98
//     16'b1111111111001110  //  -50
// };




    localparam logic signed [TWIDDLE_SIZE-1:0] TWIDDLE_REAL [0:15] = '{
        16'b01_00000000000000,
        16'b00_11111011000101,
        16'b00_11101100100001,
        16'b00_11010100110111,
        16'b00_10110101000001,
        16'b00_10001110001110,
        16'b00_01100001111110,
        16'b00_00110001111100,
        16'b00_00000000000000,
        16'b11_11001110000100,
        16'b11_10011110000010,
        16'b11_01110001110010,
        16'b11_01001010111111,
        16'b11_00101011001001,
        16'b11_00010011011111,
        16'b11_00000100111011

    };

    localparam logic signed [TWIDDLE_SIZE-1:0] TWIDDLE_IMAG [0:15] = '{
        16'b0000000000000000,
        16'b1111001110000100,
        16'b1110011110000010,
        16'b1101110001110010,
        16'b1101001010111111,
        16'b1100101011001001,
        16'b1100010011011111,
        16'b1100000100111011,
        16'b1100000000000000,
        16'b1100000100111011,
        16'b1100010011011111,
        16'b1100101011001001,
        16'b1101001010111111,
        16'b1101110001110010,
        16'b1110011110000010,
        16'b1111001110000100
    };

endpackage
